/*
 * Copyright (c) 2025 ReJ aka Renaldas Zioma
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tqvp_rejunity_vga (
    input         clk,          // Clock - the TinyQV project clock is normally set to 64MHz.
    input         rst_n,        // Reset_n - low to reset.

    input  [7:0]  ui_in,        // The input PMOD, always available.  Note that ui_in[7] is normally used for UART RX.
                                // The inputs are synchronized to the clock, note this will introduce 2 cycles of delay on the inputs.

    output [7:0]  uo_out,       // The output PMOD.  Each wire is only connected if this peripheral is selected.
                                // Note that uo_out[0] is normally used for UART TX.

    input [5:0]   address,      // Address within this peripheral's address space
    input [31:0]  data_in,      // Data in to the peripheral, bottom 8, 16 or all 32 bits are valid on write.

    // Data read and write requests from the TinyQV core.
    input [1:0]   data_write_n, // 11 = no write, 00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [1:0]   data_read_n,  // 11 = no read,  00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    
    output [31:0] data_out,     // Data out from the peripheral, bottom 8, 16 or all 32 bits are valid on read when data_ready is high.
    output        data_ready,

    output        user_interrupt  // Dedicated interrupt request for this peripheral
);
    // 256 pixel vram (16x16, ~18x14, ~25x10)
    // 256x3 = 768
    // 256x4 = 1024

    // 320 pixel vram (20x16)
    // 320x3 = 960

    // 384 pixel vram (24x16)
    // 384x2 = 768
    // 384x2.5 = 960

    // vertical
    // 192x4 = 256x3 = 384x2 = 768


    // TODO:
    assign vga_cli = (data_write_n != 2'b11); // Any write resets interrupt, TODO if need to be more careful
    // \TODO

    localparam PIXEL_COUNT      = 320;
    localparam REG_LAST_PIXEL   = PIXEL_COUNT / 8 - 1;
    localparam REG_BG_COLOR     = 6'h30;
    localparam REG_FG_COLOR     = 6'h31;
    // localparam REG_BANK         = 6'h3F;

    localparam REQ_WAIT_HBLANK  = 6'h00;
    localparam REQ_WAIT_PIXEL0  = 6'h04;
    // localparam REG_Y            = 6'h10;

    reg [PIXEL_COUNT-1:0] vram;
    reg [5:0]   bg_color;
    reg [5:0]   fg_color;

    reg         pause_cpu;
    reg         wait_hblank;
    reg         wait_pixel0;
    assign data_ready = !pause_cpu;

    always @(posedge clk) begin
        if (!rst_n) begin
            bg_color <= 6'b010000;
            fg_color <= 6'b001011;

            pause_cpu   <= 1'b0;
            wait_hblank <= 1'b0;
            wait_pixel0 <= 1'b0;
        end else begin
            // WRITE register
            if (~&data_write_n) begin
                if (address <= REG_LAST_PIXEL) begin
                    if (data_write_n == 2'b10) begin // TODO: only 32-bit writes are supported atm
                        vram[{address[5:2], 5'b00000} +: 32] <= data_in[31:0];
                    end
                end else if (address == REG_BG_COLOR) begin
                    bg_color <= data_in[5:0];
                end else if (address == REG_FG_COLOR) begin
                    fg_color <= data_in[5:0];
                end
            // READ register
            end else if (~&data_read_n) begin
                if          (address == REQ_WAIT_HBLANK) begin
                    pause_cpu   <= 1'b1;
                    wait_hblank <= 1'b1;
                    wait_pixel0 <= 1'b0;
                end else if (address == REQ_WAIT_PIXEL0) begin
                    pause_cpu   <= 1'b1;
                    wait_hblank <= 1'b0;
                    wait_pixel0 <= 1'b1;
                end
            end

            if (wait_hblank && vga_blank) begin // NOTE: do not block cpu during the VBLANK/VSYNC
                                                // TODO: block until the next blank, if already inside the blank
                pause_cpu   <= 1'b0;
                wait_hblank <= 1'b0;
            end
            if (wait_pixel0 && vram_index == 0) begin
                pause_cpu   <= 0;
                wait_pixel0 <= 0;
            end
        end
    end

    wire        vga_cli;
    wire [10:0] vga_x;
    wire  [9:0] vga_y;
    wire        vga_hsync;
    wire        vga_vsync;
    wire        vga_new_scanline;
    wire        vga_blank;

    vga_timing vga (
        .clk,
        .rst_n,
        .cli(vga_cli),
        .x(vga_x),
        .y(vga_y),
        .hsync(vga_hsync),
        .vsync(vga_vsync),
        .retrace(vga_new_scanline),
        .blank(vga_blank),
        .interrupt(user_interrupt)
    );

    reg [6:0] vga_x_per_pixel;
    reg [6:0] vga_y_per_pixel;
    reg [6:0] vram_pixel_x;
    reg [6:0] vram_pixel_y;
    reg [8:0] reset_vram_index_on_blank;

    always @(posedge clk) begin
        if (!rst_n) begin
            reset_vram_index_on_blank 
                            <= 9'd0;
            vram_index      <= 9'd0;
            vram_pixel_x    <= 7'd0;
            vram_pixel_y    <= 7'd0;
            vga_x_per_pixel <= 7'd57 - 1; // 1024/18=~56  (18x14 = 252)
            // vga_y_per_pixel <= 7'd56 - 1; // 768/14 =~56
            // vga_y_per_pixel <= 7'd4 - 1;
            vga_y_per_pixel <= 7'd2 - 1;
        end else if (vga_new_scanline) begin
            vram_pixel_x <= 7'd0;
            vram_index   <= reset_vram_index_on_blank;
            if (vram_pixel_y == vga_y_per_pixel) begin
                if (vram_index == PIXEL_COUNT-1) begin
                    reset_vram_index_on_blank <= 9'd0;
                end else begin
                    reset_vram_index_on_blank <= vram_index + 9'd1;
                end
                vram_pixel_y <= 7'd0;
            end else begin
                vram_pixel_y <= vram_pixel_y + 7'd1;
            end
        end else if (vga_blank) begin
            vram_pixel_x <= 7'd0;
        end else begin
            if (vram_pixel_x == vga_x_per_pixel) begin
                vram_index   <= vram_index + 9'd1;
                vram_pixel_x <= 7'd0;
            end else begin
                vram_pixel_x <= vram_pixel_x + 7'd1;
            end

            if (vram_index == PIXEL_COUNT-1) begin
                vram_index   <= 9'd0;
            end
        end
    end

    reg [8:0] vram_index;
    // always @(posedge clk) begin
    //     if (!rst_n) begin
    //         vram_index <= 9'd0;
    //     end else if (vram_index == PIXEL_COUNT-1) begin
    //         vram_index <= 9'd0;
    //     end else begin
    //         vram_index <= vram_index + 9'd1;
    //     end
    // end


    reg pixel;
    reg hsync_buf;
    reg vsync_buf;

    always @(posedge clk) begin
        if (!rst_n) begin
            pixel <= 1'b0;
        end else if (vga_blank) begin
            pixel <= 1'b0;
        end else begin
            pixel <= vram[vram_index];
        end
        hsync_buf <= vga_hsync;
        vsync_buf <= vga_vsync;
    end


    wire [5:0] rrggbb = pixel ? fg_color : bg_color;
    assign uo_out = {hsync_buf, rrggbb[5:3], vsync_buf, rrggbb[2:0]};
    assign data_out = {22'd0, vga_y};

    // List all unused inputs to prevent warnings
    wire _unused = &{ui_in, 1'b0};

endmodule
